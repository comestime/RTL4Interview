../Mem_Access/FIFO_1Port_RAM.sv