../FIFO/fifo_async_even_entry.sv