../Mem_Access/FIFO_Dual_Port_RAM.sv